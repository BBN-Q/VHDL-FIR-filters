package DataTypes is
  type integer_vector is array(natural range <>) of integer;
end DataTypes;
