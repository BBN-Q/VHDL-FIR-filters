package DataTypes is

  --VHDL 2008 compatibility definitions
  type integer_vector is array (natural range <>) of integer;
	type real_vector is array (natural range <>) of real;

end DataTypes;
