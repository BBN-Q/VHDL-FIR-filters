library ieee_proposed;
use ieee_proposed.standard_additions.all;

package TestVectors is

--Generated in Julia with
-- freqs = [linspace(0,0.49,1024); linspace(0.49,0,1024)]
-- phases = cumsum(2pi*freqs)
-- chirp = sin(phases)
-- writecsv("chirp.dat", reshape(chirp, 16, 128)')

--Then add leading zeros to numbers

constant chirp : real_vector(0 to 2047) := (0.0,0.003009536806409242,0.00902850138597494,0.01805626680915896,0.030090870627762445,0.04512778893385701,0.06315830334398528,0.08416746365467088,0.1081316513467636,0.13501575270392485,0.1647699552745627,0.19732618795505588,0.23259423329540294,0.27045755089024237,0.3107688630451513,0.35334556837680536,
0.3979650656271231,0.44436008867398213,0.492214174329677,0.541157406733794,0.5907626055234261,0.6405421488846443,0.6899456462472261,0.7383586977611637,0.7851029975439158,0.8294380535330721,0.8705648069085382,0.9076314365305237,0.9397416265532694,0.9659655560560904,0.985353835847693,0.9969545672357113,
0.9998336283478008,0.993098203681623,0.9759234605714718,0.9475821415081322,0.9074766839868438,0.8551733012222782,0.7904372605414078,0.7132683861265141,0.6239355955404599,0.5230090637416955,0.41138840491780465,0.29032508447857214,0.16143713607489332,0.026714178440184432,-0.11148927766353814,-0.2504741524056887,
-0.38723246764555697,-0.5184997523888724,-0.6408250967390806,-0.750659144632319,-0.844459540256473,-0.9188124230713243,-0.9705675197106018,-0.9969832380393471,-0.9958769731678246,-0.9657746454868569,-0.906052379102604,-0.8170622805683274,-0.7002335879567966,-0.5581401307030633,-0.3945251734097812,-0.21427540733029884,
-0.023337181410284943,0.17142991496745547,0.36246427460134084,0.5417770443832358,0.7012851793704834,0.8331930511332957,0.9304081884205805,0.9869720849674907,0.998482762710716,0.9624823231047318,0.878780476678668,0.7496844325171813,0.5801069390895341,0.37752800094067573,0.15179203288285922,-0.08526903490336298,
-0.32038512175441497,-0.5395553163566308,-0.7288845332352496,-0.8755065743515619,-0.9685373216766484,-0.9999907578314463,-0.9655832102953302,-0.8653490020710597,-0.7039947321236275,-0.49093050801619365,-0.2399348967121132,0.03156423096859243,0.3035795606948041,0.554976423542041,0.76512246825717,0.9156564214027707,
0.992229748283805,0.9860574269475277,0.8951101416022761,0.7247927872291202,0.4879847538944498,0.2043657872951862,-0.10098500800378113,-0.3996547696896962,-0.6624858701313991,-0.8624722260556263,-0.9776854982698263,-0.9939153764222104,-0.9067010731116909,-0.7224612869978785,-0.45849945797668906,-0.14176767008861546,
0.19359164833596,0.5097549329851089,0.7694551316729513,0.940495268869067,0.9999971311523873,0.9378161098720055,0.7585980726597946,0.4820765737729079,0.14140286722282824,-0.22045032082258614,-0.5558957502485246,-0.8189699885509141,-0.9718115683235424,-0.9904665028066892,-0.8691103911628966,-0.6219176215726087,
-0.28208612551292306,0.10208484025991485,0.47371412522620115,0.7756556741932306,0.9594410459527343,0.9934537003170656,0.8689280578080635,0.6025913882102425,0.2352217084180098,-0.17397076096020336,-0.556508257325929,-0.846034939448263,-0.9900819874211214,-0.960113564153681,-0.757877281039339,-0.41658791360854364,
0.0036851443318938774,0.42600157376882175,0.7703957794606774,0.9691760809730396,0.9807598096756696,0.7991588502212595,0.4568611927796644,0.020021325011503454,-0.42361069535174145,-0.7820119797363023,-0.9781476007338062,-0.9671468547019576,-0.747485377619804,-0.3632655363652322,0.10355108894709533,0.5499080320410813,
0.8741975405992937,0.999747348223655,0.8937918478707404,0.57710130140866,0.12131051127045517,-0.36623929527092397,-0.7672537884830104,-0.9813074417843966,-0.9517374557985222,-0.6818111745341409,-0.23635577000374525,0.27252648258092055,0.712923914654375,0.9672872319411949,0.9645209437798339,0.7011100198920515,
0.2447615401491162,-0.28155575815508593,-0.731904985133538,-0.977827203469026,-0.9458014962845844,-0.6406364745033382,-0.14705512309060723,0.3923229928796036,0.8174162385389457,0.9983691039261356,0.8763066800438617,0.48412008290905373,-0.060399719116204925,-0.5885303405240491,-0.9324200145421188,-0.9790449513348892,
-0.7088635043456892,-0.20556809148195004,0.36795322802146924,0.8212893954598222,0.999851070636544,0.8388545022400569,0.38876087467720755,-0.19828947779701137,-0.7184147473419972,-0.9865236332696655,-0.9032254930442208,-0.49365702039443676,0.09750139798951075,0.6553247858262308,0.9722299502635644,0.9261372306899166,
0.529537243230223,-0.07087970523087107,-0.6464657272875212,-0.9730149601055464,-0.9190304590967838,-0.5008508079896566,0.11917643640146519,0.6936267608545286,0.9881310876402234,0.8781348357467017,0.4039854524222203,-0.24082917116248592,-0.7866222636324429,-0.9999999320982497,-0.7852171069867128,-0.2298455115386206,
0.42794544478660324,0.8998236566283769,0.9739562425374275,0.6122516786220964,-0.027266749953944257,-0.6567154575126752,-0.9868829976729444,-0.8612574561354325,-0.33303962284887434,0.3538626294741027,0.8752393373095374,0.9795917130443866,0.6116687696549368,-0.055065166571763094,-0.6971137303000885,-0.9967895420987216,
-0.8008172096917993,-0.2019602556167706,0.5011697363315456,0.950942574239053,0.913170348342943,0.4019618364271304,-0.32090870757079654,-0.8772223479476128,-0.9699878658804659,-0.5445102523831808,0.1756640161845937,0.8027991649817908,0.9928584451589106,0.6363822732171698,-0.07455509966342397,-0.7460147715278668,
-0.9991305290471304,-0.6857550264239899,0.020819608243733,0.7175597230268717,0.9999282796327078,0.6985215078380845,-0.015169963271232486,-0.7219939967957573,-0.9995378793034809,-0.6764011186838979,0.057640673498476395,0.758638089460936,0.9953010338365573,0.616467802601186,-0.14778410084196264,-0.8214295322152841,
-0.9776725938491636,-0.5119725209679009,0.2832055066823071,0.8978045395707454,0.9306556045244803,0.3546667317622784,-0.4565333534321916,-0.9671468547019587,-0.8333628305021649,-0.139031182736121,0.6512326646894941,0.9999511092514303,0.6638649715342271,-0.13136343479314716,-0.8373803493776546,-0.9595448687006312,
-0.4065121938376615,0.4359774574035154,0.9696734391395803,0.8086919590317078,0.06309700663582171,-0.7302287195504364,-0.9912128323494174,-0.5229567134958419,0.3339660692878813,0.9439311361895816,0.8470484776098806,0.11032951228390593,-0.7119757308619643,-0.9918976940185701,-0.5094378574515116,0.36846716451084466,
0.9614589591440175,0.8024694517660159,0.010502492033069953,-0.791602106251714,-0.9638857899292189,-0.36280770535064155,0.5326077245748038,0.9973257110483206,0.6480107572161985,-0.23480381542571258,-0.9253708340230731,-0.8476681608676327,-0.06052233281288099,0.7792481574010718,0.9611374492925813,0.325035767005935,
-0.5907626055234363,-0.9996281930532712,-0.5433764119924255,0.3872324676455613,0.9804468152472404,0.7108966714680653,-0.1891909347174483,-0.9224807993526507,-0.8305001189027361,0.010133996385618384,0.8432401600228956,0.9095299100544573,0.14249721801298765,-0.7573160248834863,-0.9572129199008955,-0.2657830970450335,
0.6759033540093659,0.9828240714433278,0.35971506046498386,-0.6069935629405327,-0.994521895368272,-0.4257792915650477,0.5558957502485402,0.9987040337033605,0.46585230769898595,-0.5258330419974852,-0.9997072143929236,-0.4814307090066736,0.5184472332082753,0.9996982296182911,0.4731731300150035,-0.5341143830265777,
-0.9986471571584262,-0.44072497632647023,0.5720241321969255,0.9943276055603799,0.38281110260288054,-0.6300122509251622,-0.9823447484717093,-0.29760454137079934,0.7041691918475176,0.9562478732841506,0.18339791961086335,-0.7882879722427368,-0.9078375815147489,-0.039605030117346514,0.8732714326171994,0.8278220913767712,
-0.13191139741955799,-0.9466954347721885,-0.7069981979993822,0.32526809421017217,0.9928144144618846,0.5381065856032361,-0.5289640103269578,-0.9933762948065417,-0.31840624874680734,0.7246658275120037,0.929640763239943,0.0527959634614048,-0.8869990161229342,-0.7859012036730183,0.24303417259179474,0.9851330761850796,
0.5545165057524383,-0.5403824463241964,-0.9869424227098641,-0.24190203061626359,0.7976425852718727,0.8661789109735056,-0.12588162850958684,-0.9643423579907037,-0.6122516786220984,0.5002127472973367,0.9903817087026202,0.24082917116249067,-0.8125760460551121,-0.8405222389558581,0.19822927778232555,0.9855105177336685,
0.511919760787658,-0.6205218425053521,-0.9528060927220973,-0.0494836673941917,0.9193207369594582,0.6862912748432994,-0.44886626208371305,-0.9928584451589092,-0.22146863967111008,0.8455434164577524,0.7833881594814794,-0.33049023947582035,-0.9999822531753753,-0.31636772331629964,0.7980498849413383,0.8240827009128945,
-0.27961034302780163,-0.9994742149208529,-0.33842006607345415,0.7930260663301479,0.8202367903138472,-0.300476366013053,-0.9999902221637745,-0.2891493903803436,0.8320023962994877,0.7706306799313083,-0.39147540029082745,-0.9932201235392927,-0.1654362947032718,0.9022213898145305,0.6613349006269055,-0.5434279717304601,
-0.9541944001434448,0.03616802537012879,0.9740119169423311,0.4707364456244408,-0.7325324463663174,-0.8438339163645456,0.3086664945538131,0.9979409733823245,0.1814050879186457,-0.9106244488419474,-0.6183038120094322,0.6183520826077329,0.9080949545204179,-0.19919238812883314,-0.9996078251217901,-0.2508309036018743,
0.8888073030669474,0.6408250967390567,-0.6121059825476693,-0.9025125569326886,0.23259423329540876,0.9996281930532709,0.17626862454778633,-0.9291647398852818,-0.5455916271926222,0.7161465663659762,0.8220245602068306,-0.40449104820502535,-0.9736629875454723,0.046600298701223,0.9910659887014124,0.3061533553493653,
-0.8844329309978163,-0.6106478796354173,0.6783890876748908,0.8363380688609343,-0.40583869896206176,-0.9667553674955928,0.10208484025992764,0.9986977743648844,0.1999747736860411,-0.9398465739188324,-0.47317313001499317,0.8055736181852027,0.6978619477542214,-0.6155969412627498,-0.8623478618976288,0.39096668520026323,
0.962298780113776,-0.15167061671144172,-0.9994860956681558,-0.08502425025169756,0.9802043489236637,0.30551011556746877,-0.9136453558472694,-0.500159563302943,0.8104226230378767,0.6631757022752622,-0.6813617471053987,-0.7921272252122072,0.5366044367994838,0.8873107915913352,-0.3850228896961935,-0.9510565162951624,
0.23390818439176708,0.9870608706849536,-0.08887900284181341,-0.9998007809911357,-0.04604811923255608,0.9940566168239611,0.16828252699735496,-0.9745516609908547,-0.27642446243820146,0.9457017236776248,0.37000829782270866,-0.9114601364290008,-0.44925040958431006,0.8752393373095212,0.5148186974659404,-0.839889431929051,
-0.5676330748505911,0.8077153707864679,0.6087005182942585,-0.7805168041851936,-0.6389843818080108,0.759637579003864,0.6593054089160205,-0.7460147715278446,-0.6702709013310781,0.7402198481609974,0.6722285105447275,-0.74248690716596,-0.6652418190580283,0.7527249895692291,0.6490860223763096,-0.7705132427757734,
-0.6232633982105118,0.7950794082574641,0.5870396651653683,-0.8252638349728042,-0.5395036034246844,0.8594731360198571,0.4796532334934171,-0.8956298176088092,-0.4065121938377049,0.9311267646589968,0.31927945262819196,-0.9627983170842194,-0.21751382568137756,0.9869226292560654,0.10135163253635993,-0.9992727076427971,
0.0282490786318487,0.995235387930964,-0.16925113838257813,-0.9700177271331867,0.3182898011272373,0.918957811620246,-0.4704654806027301,-0.8379506339882749,0.6192205543224406,0.723988293607887,-0.7563525689854483,-0.5757964221204458,0.8722220221371341,0.3945251734098272,-0.9562119287439873,-0.18442423636280345,
0.9974848707556324,-0.046600298701206355,-0.986057426947534,0.2866790147178757,0.9141689165592279,-0.5200744174014562,-0.7778605283231228,0.727832428333732,0.5786051024563174,-0.8891167201038921,-0.3247453304142152,0.9832856736347091,0.03242365970004785,-0.9926592452937683,0.2743579135376505,0.9057662769001549,
-0.5648994311036025,-0.7206753156820325,0.8044440495242888,0.44782315797847155,-0.9583605839469564,-0.11161134942519921,0.9976264831905004,-0.249998431239785,-0.9049838971925831,0.5885303405239972,0.6807321169304228,-0.8509751277299115,-0.3467868358438891,0.9884217748453573,-0.052489293221122,-0.9662983868680873,
0.4539631370664746,0.7743748328218639,-0.7845320505833934,-0.434041837571043,0.9745516609908637,0.00018425763267310779,-0.9739562425374421,0.44452514801095727,0.7676869123472986,-0.803713747636311,-0.3860429701803985,0.9884124537627461,-0.09444461441083994,-0.9412235685085133,0.5626166466134139,0.6573173897703839,
-0.8968285939042069,-0.19497737248848954,0.9976349340503157,-0.3304902394757889,-0.8208686878033611,0.771959804857379,0.4002739881798558,-0.9913342766188038,0.150759922603009,0.9058443457811144,-0.6642782626614976,-0.5245263618332162,0.9671468547019388,-0.04107789109591492,-0.9420093690481555,0.6022972537332242,
0.5788054609516353,-0.9532154263569601,0.006080464441631211,0.9485199833983428,-0.598367660536584,-0.5705118131163525,0.9605246836315129,-0.046293534076723965,-0.9295728545714914,0.6531881029862465,0.498403434215545,-0.983575166388413,0.16107344366955956,0.87369006714982,-0.7561114481407832,-0.35334556837688336,
0.9999829774565238,-0.34523094969406093,-0.7558702246135975,0.8810856808552074,0.12496761564785265,-0.9701221262494077,0.579756686516427,0.5446647900005732,-0.9807358219647636,0.18472605601723924,0.8412535328311919,-0.8189699885509125,-0.21799338873123264,0.9847828571196285,-0.5414156248318981,-0.5631750581513363,
0.9810940835735036,-0.21013400304633442,-0.8131841776087743,0.8591904377672706,0.12131051127042962,-0.9562478732841403,0.6581963830082829,0.41491212964399315,-0.9999999528460065,0.417090373258072,0.6495531250812842,-0.9636564368049945,0.16834306997976228,0.8186526622612009,-0.8710479313477645,-0.0648132236470992,
0.9261372306899257,-0.74556469186207,-0.2684465346908975,0.9822181311559998,-0.6071887856666901,-0.4364196022375329,0.9998369723254462,-0.4712782424595576,-0.5682397043447859,0.9921147013144757,-0.34857204732177216,-0.6668910543849532,0.9707889808499951,-0.24589284302943243,-0.7369902686188161,0.9454418975268769,
-0.16713208997710216,-0.7833881594814752,0.9232613490220778,-0.11423548190615558,-0.8102066749327611,0.9090954351636021,-0.08802250412435592,-0.8202367903138108,0.9056100468861878,-0.0887566498907658,-0.8146115771517082,0.9134205073483317,-0.11643181800740429,-0.7926892027355031,0.9311267646590053,-0.17076426610548007,
-0.752118153880495,0.9552359739505435,-0.250890358824081,-0.6891004559833478,0.9800093109258199,-0.35478158212489985,-0.5989088383564629,0.9973257110483137,-0.47841322123045255,-0.4767403902519586,0.9967153549717618,-0.6147737702287474,-0.3189884147417508,0.9657746454868743,-0.7528867045390852,-0.12496761564792558,
0.8912155576862733,-0.8771338738564847,0.10098500800376188,0.760794742955482,-0.9673028111683966,0.34730525284481817,0.5662670316000387,-0.9998849294865633,0.5934353651266506,0.307264076565365,-0.9511513693477767,0.809341782516656,-0.004422168794159757,-0.8023228338466111,0.9573904770607453,-0.3412504929989564,
-0.5466206641503774,0.9976264831904988,-0.6587510748834505,-0.19708533568323386,0.8969915561254791,-0.8988568606925815,0.20713062292343057,0.6418147286455205,-0.9995921928281882,0.5994005809751299,0.2510092664292314,-0.9116116774438707,0.8929916135407523,-0.21481530836810034,-0.6193652260561446,0.999770272652233,
-0.6547214702012885,-0.16089158926103178,0.8593475247690308,-0.9452015230229605,0.36332275907767175,0.4719823125318807,-0.9761373308268763,0.8030188375198256,-0.07792332300584576,-0.6985215078381339,0.9987071577214577,-0.6246073315482653,-0.16688986365536693,0.8452153357308497,-0.963112999918026,0.44848203161303646,
0.35713483232269194,-0.9292782190132033,0.9022213898145017,-0.29901148777082964,-0.4921607095671134,0.9710976421195604,-0.8412535328311632,0.1892512443603208,0.577602786377844,-0.9884962092722293,0.7970865899203154,-0.12496761564780015,-0.6200882692064322,0.9938679288387599,-0.7792481574010551,0.10813165134672571,
0.6239355955405227,-0.993054914643193,0.7911139717062325,-0.13909200518191323,-0.5895726246997116,0.9850379631877175,-0.8304659057025278,0.2171541189252232,0.5133963151420596,-0.961980716781132,0.8891167201038432,-0.33951794380192696,-0.3890437958192758,0.9097085232999785,-0.9517939907728709,0.49866964616791687,
0.2103141431167259,-0.8092335472757787,0.9950051160607164,-0.6786146800234728,0.02395120180730649,0.6403534686527573,-0.9872375372801687,0.850975127729915,-0.3031113592779437,-0.3884213209136557,0.8924657858207963,-0.973014960105543,0.5972844857682161,0.05469720669896284,-0.6791107578847878,0.9908434520759539,
-0.8523271198571188,0.33124371843148886,0.3355287158596355,-0.8515552468448278,0.9925773071348301,-0.7019416503485776,0.11014637765939872,0.5264075886970603,-0.9377521321470998,0.9541392564000708,-0.5737357457973932,-0.04163019112336702,0.637565951874243,-0.9730291302641741,0.9167638907170019,-0.4962187255104266,
-0.11813968643030039,0.6838752253402491,-0.9827332759560277,0.9036731045547635,-0.48175367410166126,-0.11966427385297947,0.6739545885325248,-0.9770488453596863,0.9214818920953487,-0.5322957910160776,-0.04623218062730768,0.6058214576322056,-0.9497191599602935,0.9610356479162242,-0.640542148884525,0.10251251918187369,
0.4678076793701199,-0.878780476678683,0.9963054041344797,-0.7860151264228127,0.3210832143937779,0.24505928381262787,-0.7304804406102583,0.9832409137134386,-0.9278877894237486,0.5861443029616399,-0.06683566150860297,-0.47019447121243707,0.8638677340617551,-0.9997473482236539,0.8419832907437576,-0.4408903662690388,
-0.0846570636566797,0.5835536806699074,-0.9161741113769784,0.9928144144618726,-0.7965299180241628,0.3850228896961691,0.1277093329230095,-0.6038650247938312,0.9190304590968579,-0.9940566168239582,0.813684326191554,-0.4279454447865235,-0.06297441250568013,0.5356193469900112,-0.8745253979533913,0.9999486497402055,
-0.8855767543105344,0.5626166466134528,-0.11014637765932567,-0.3651531610394594,0.7545416612274612,-0.971883923136893,0.9719417409952203,-0.758638089460823,0.38213011024830146,0.07394260288837638,-0.5116559309237626,0.8399560970716563,-0.9932201235393043,0.9435655718586581,-0.7048230371960105,0.32793844246439097,
0.11069577028933286,-0.5252059900505713,0.837111664224536,-0.9898214418809346,0.9581850139827753,-0.7516727352889859,0.4110524900156274,0.0003685152590503231,-0.4089797830029079,0.7441713858688352,-0.950313584945024,0.9954543908729976,-0.8755065743514975,0.6135620073069442,-0.25481230017595263,-0.14176767008867705,
0.5133963151421858,-0.8034212872505613,0.9696734391395753,-0.9900819874211002,0.8649177419171217,-0.6155969412626711,0.28049476550663527,0.09138694014486592,-0.44782315797844435,0.740715200538672,-0.9323756165982682,0.9999815138052176,-0.9377521321470722,0.7567542087874055,-0.4825608005139252,0.15124564210050895,
0.19563997275486703,-0.5163974616389775,0.774141610639138,-0.9408287453232455,0.9999592422507653,-0.9477586144480888,0.7928389497974999,-0.554516505752347,0.2600943367236547,0.058499091417676743,-0.3682958648498571,0.6387008692197899,-0.844393739249907,0.9674739418226755,-0.998707157721458,0.9378374287048756,
-0.793026066330077,0.5795564940700957,-0.31799866106999747,0.03205533599918914,0.25368368280914405,-0.5158714014515795,0.7342443331796533,-0.8930468930979533,0.981963551580303,-0.9965338543740583,0.938071702353161,-0.8131484296986246,0.6327271278299932,-0.411052490015664,0.1644064656851177,0.09016362750488506,
-0.3360493932155833,0.5581401307031082,-0.743678855697571,0.8828803031216433,-0.9692970183318317,0.9999388890464364,-0.9751674941476394,0.8983987903338475,-0.7756556741931248,0.6150159489703182,-0.42600157376871184,0.21895235682583444,-0.004422168794093122,-0.20737096559408913,0.4070171700992913,-0.5862935797755201,
0.7384415354309304,-0.8583407681610312,0.9425850967230406,-0.989468820491541,0.9988963752162109,-0.9722299502635492,0.9120907404896746,-0.8221294721367157,0.7067809816208303,-0.5710161349452881,0.4201024494335945,-0.25938260183508033,0.09407773995878312,0.07087970523103725,-0.23098107678529725,0.38224362339952933,
-0.521280465089599,0.6453404007414902,-0.7523205033996403,0.8407550898971677,-0.9097850203600489,0.9591114143970019,-0.9889378035353178,0.9999045146821158,-0.9930187374259302,0.9695833066135923,-0.9311267646589543,0.8793367845001981,-0.815998557859173,0.7429393030681001,-0.6619796358202397,0.5748921838049382,
-0.48336751734237515,0.3889872145252193,-0.29320367996313995,0.19732618795504092,-0.10251251918199361,0.009765499361732759,0.08006627731206205,-0.16628425381335468,0.2483329326039654,-0.3257907586179394,0.39835945097007797,-0.4658523076990683,0.5281819400392355,-0.585347823987661,0.6374239897487832,-0.6845471059287667,
0.7289686274213192,-0.7724281043368765,0.8142908406281377,-0.8538653082573495,0.8904062471387754,-0.9231197129162523,0.9511703291944407,-0.973690986386355,0.9897952024830696,-0.9985923196736443,0.9992056528127146,-0.9907936294308838,0.9725738648749349,-0.9438499993586177,0.9040409860797071,-0.8527123619742235,
0.7896088572172193,-0.7146875097917164,0.6281502525425606,-0.5304747392193905,0.4224419821687822,-0.30515919870949115,0.1800761189395576,-0.048992909692217416,-0.08594216611389639,0.22224719123044084,-0.35713483232250426,0.4875558158792575,-0.6102587018467122,0.7218664968088648,-0.8189699885508276,0.8982368845725034,
-0.9565349101126893,0.9910659887013882,-0.9995075245064499,0.980155678160314,-0.9320644370998785,0.8551733012223655,-0.7504156194341595,0.619799115069694,-0.4664500244525497,0.29461263699310736,-0.10959695137365037,-0.08233128363368569,0.27412165561340135,-0.45817192929087336,0.6266197666740837,-0.7716864364913274,
0.8860612610601908,-0.963311071228459,0.9982946401623997,-0.9875582919900078,0.929686018151282,-0.825575885921291,0.6786146800236204,-0.49472492022941666,0.2822628954861536,-0.05175326450312388,-0.18454496631315256,0.4132349370166846,-0.6205218425051876,0.7930634806625457,-0.9188851329441853,0.9883003099499879,
-0.9947694241718418,0.9356230194382439,-0.8125760460552138,0.6319658385734424,-0.4046595526747851,0.14559692833675505,0.12703922465371412,-0.3930008272302543,0.6314420981441912,-0.8225837679155386,0.9494495813049737,-0.9995266093703139,0.9661876218509289,-0.8497146358473731,0.6577801294488398,-0.4052772848121739,
0.11344222272220064,0.19172332242894882,-0.48164602633714915,0.7278324283337864,-0.9047485840218507,0.9926443811472276,-0.9800093109258532,0.8653490020711206,-0.6580114062480836,0.37786921976079496,-0.0537772746282929,-0.27913855395156517,0.5831545944078496,-0.8222343561547691,0.9664563127610382,-0.996042430247767,
0.904434403102149,-0.6999265870895341,0.40550186882994016,-0.0567208927375932,-0.3022332844683147,0.6239835919886342,-0.8642387554651628,0.988112210606618,-0.9755739114024538,0.825159761948515,-0.5552318601600674,0.20238131206587956,0.18303564237474998,-0.5437888324861159,0.8242218444828765,-0.9790449513348735,
0.981082195177678,-0.8266142333279635,0.5372262223602278,-0.15755663003235412,-0.2510092664289591,0.6199437026616289,-0.8850626948616677,0.9980035213959386,-0.9356230194381778,0.7054327531260632,-0.345749684110091,-0.07988260987170116,0.4933899289830585,-0.8163179657269587,0.984942549204219,-0.9634263711776858,
0.7522395721049543,-0.38977921901305135,-0.05365461355289506,0.4888422763808734,-0.8253678799787844,0.990651734593477,-0.9462791630151721,0.6978619477543273,-0.29578627897704307,-0.17397076096015773,0.6075791211626508,-0.9061822888493543,0.9988702597427269,-0.8604135663527708,0.5191823236734671,-0.052673295961159876,
-0.42911081873596063,0.809161375184775,-0.9920915908679907,0.928892032477951,-0.6312515756066563,0.1710668434510288,0.3357022863775637,-0.7575967229797923,0.9818355894364744,-0.9452616647897176,0.6534206039901576,-0.18176747662336665,-0.3424625884345986,0.7738304841968899,-0.9891282984389744,0.9234735680832437,
-0.5913075845621006,0.08520783922241884,0.4484820316130653,-0.851297544578493,0.9999917838993665,-0.8454122224360152,0.43038636152649234,0.12021305644662868,-0.6357187576162566,0.9522075930817174,-0.9653431787143063,0.6663416711426023,-0.14827004143491054,-0.42110544953640666,0.852712361974076,-0.9992056528127103,
0.8066276677025832,-0.33622292952380883,-0.2528518488647115,0.7559908492104458,-0.9940566168239405,0.8783110786918841,-0.4455151869048634,-0.15124564210075886,0.6949970166042289,-0.9833415400775091,0.9048270524661484,-0.48412008290920405,-0.1229564150817109,0.6852184054929852,-0.983619481132019,0.8976421866433947,
-0.4562054520857639,-0.16913007087895782,0.7288424820177626,-0.9945475455778356,0.8534494477966422,-0.35868329784557457,-0.2877379816955846,0.8155012056206679,-0.9988702597427072,0.7549043043342549,-0.18369979828393643,-0.46976076396498595,0.9191030753715493,-0.9624823231047431,0.5754950874891336,0.07253375482952198,
-0.6899456462474445,0.993098203681613,-0.8379506339882754,0.2913828346595179,0.39418652342810256,-0.8952743815374141,0.9701072230683514,-0.577602786377572,-0.09695124396905688,0.726356599131414,-0.999244331726306,0.7756556741931081,-0.16210384850817697,-0.5355156108715252,0.9624989870476973,-0.8963934326111725,
0.36589635932450076,0.35730693262553836,-0.8949731821311325,0.9600620275154005,-0.5126054924302825,-0.2121751712905391,0.8242218444829597,-0.9878463667270956,0.6081155929384682,0.11014637765935094,-0.769101957602283,0.9970590315798641,-0.6601362383507253,-0.05506516657171462,0.7407564617448984,-0.9989645242676494,
0.6744082097959153,0.047950010449071295,-0.7440482912135733,0.9980497999250735,-0.6527229161979853,-0.08887900284209549,0.778439169653416,-0.9918742692338919,0.5923967326822825,0.17723585952633023,-0.8378835890844295,0.9711416047200888,-0.4870731199174164,-0.3103018009850331,0.9097850203599656,-0.920188573590739,
0.32904064971048963,0.48029981659468185,-0.9735508452672408,0.8186173883419711,-0.11344222272232042,-0.6703164802773574,0.9998849294865668,-0.6451996362786244,-0.15543344474071766,0.8502323509264288,-0.9526381366075729,0.38519293582369607,0.4564240598699014,-0.9749220545325264,0.7954889886484294,-0.04138472600501908,
-0.7446635117954294,0.988215849773712,-0.5052565935761911,-0.3530008009869042,0.9503135849449365,-0.8365063837916014,0.0912646150556396,0.7250466328368242,-0.9893886575662012,0.49381725289623984,0.3848528304968512,-0.966076678240067,0.7922396745191796,0.006080464441436143,-0.8014053750519418,0.9595448687006682,
-0.3483417683229027,-0.5453342392583306,0.9982946401624035,-0.6369979735451349,-0.2483924273738288,0.9304532047581092,-0.8405555128891873,0.047643265378157953,0.7870392298417999,-0.9577091697847773,0.3138612488009501,0.5999412366881157,-0.9992656645523615,0.5343739805961967,0.39672509027439745,-0.9823562369032812,
0.7041255809007728,0.19822927778224098,-0.9258589810318574,0.8257491385636337,0.018240494096170616,-0.8473747705366452,0.9064418519499452,-0.1355634434579283,-0.761631182746552,0.9553812231416792,-0.26009433672370674,-0.6799668893964009,0.9818588886167654,-0.3552409300243176,-0.6105019552361243,0.994090001756381,
-0.4224419821685521,-0.5586496492780302,0.9985496505565259,-0.46356816289332564,-0.5277124826373812,0.9996609329070537,-0.4801381952657299,-0.5193922790374974,0.9996798527827121,-0.4728484471973341,-0.5341143830263365,0.9986662516299646,-0.4413864462632654,-0.5711169734685645,0.9944833075048162,-0.3845126729060184,
-0.6282936112808929,0.9828240714433175,-0.30041778446244793,-0.70181040379821,0.9573194975321502,-0.18738131458586693,-0.7855592753467591,0.9098360012401582,-0.04475964604561805,-0.8705648069084067,0.8311154206536021,0.12569883445977326,-0.9445378460715312,0.7119326006987798,0.31828980112732186,-0.9918586340023885,
0.5449223116007818,0.5217521137593025,-0.9943537059304711,0.3271260039055301,0.7180301204725409,-0.9332609015006821,0.06309700663579436,0.8820135345469781,-0.7926892027356017,-0.23193709834561324,0.983038759705054,-0.5645953087828166,-0.5297977237530118,0.9889378035353379,-0.25475290789969895,-0.7893449719353189,
0.873091820144023,0.11161134942490603,-0.9603365128905524,0.6241275672095501,0.48675123991752783,-0.9924497843002607,0.25653425714528477,0.8027991649816546,-0.849585078842166,-0.18122388432475217,0.9823562369033162,-0.5273472376157543,-0.6059680428363621,0.9583430432180865,-0.06861272900334009,-0.9114601364290141,
0.7006281131612322,0.4306635398763881,-0.9951088024945819,0.24190203061622081,0.8339394923866496,-0.7967155504654506,-0.3095426654061482,0.9998635186987476,-0.3379576638045487,-0.7838460353002926,0.8372124448443048,0.25653425714510186,-0.9983900742330467,0.3615482187460764,0.7775130265849035,-0.834515245110074,
-0.27577511283482764,0.9997636433157151,-0.3144443458495692,-0.8167788922655665,0.7877207631984187,0.3658963593248227,-0.9960859810354937,0.19335061331790343,0.8894538031009853,-0.6828887506604517,-0.5184472332083373,0.9626986711387306,0.0059576282447293795,-0.9666296101531855,0.49781760250371404,0.7108534742129297,
-0.8604135663526209,-0.2780177850102128,0.9994958926054978,-0.2135554374603414,-0.8964206555574948,0.6443076195263534,0.5913571147310979,-0.921910746436548,-0.16513342248771476,0.9980151418538545,-0.28491329175442515,-0.8718612961488524,0.6681258416964581,0.5828551873129414,-0.9177668215062932,-0.19624225914961008,
0.9999467654994565,-0.21349543472967644,-0.9143182260406801,0.5776027863778561,0.6883434376322585,-0.8438339163646503,-0.3677818908658628,0.9820331601986976,0.006080464441810514,-0.9847828571196761,0.345173306022015,0.8642387554650618,-0.6433677066385753,-0.6466531452122254,0.8590018264087934,0.3660678335121018,
-0.9769571724038557,-0.05837646291988922,0.9954660824282814,-0.2434511941829606,-0.9235442450681245,0.5126054924305813,0.7776675011386273,-0.7301028218305842,-0.578354605228324,0.8850912821049326,0.34713245896123557,-0.9741369694026344,-0.10416195967625463,0.9998685450900184,-0.13337243358077683,-0.9693272161076925,
0.35213867288246026,0.8922994824279628,-0.5429122821330804,-0.7798252121859228,0.700365120137631,0.642991469581631,-0.8225488407010535,-0.4920537744723097,0.9102179201840287,0.33587584549828825,-0.9661083946372618,-0.18164668312879856,0.9942555200963364,0.03481765419041372,-0.9994022053984573,0.1008016905915291,
0.9865236332696867,-0.22284598065690758,-0.9604734078158236,0.3301424088658707,0.9257428952286811,-0.42244198216862494,-0.8863173735938427,0.5001595633030974,0.8456089943312611,-0.5641389815502341,-0.8064461175055057,0.6154517245273631,0.7711001668778155,-0.6552319952211744,-0.7413338251508339,0.6845471059287581,
0.718457470112557,-0.7043000087492173,-0.7033837885419907,0.7151598988617396,0.6966732473191903,-0.7175169433783835,-0.6985654574360785,0.7114579916885062,0.7089934576382542,-0.6967613649452509,-0.7275796677215648,0.6729102950772814,0.7536138594172214,-0.6391261055633592,-0.786015126422754,0.5944236210714182,
0.8232816603908748,-0.5376923700363918,-0.8634342826731501,0.46780767937020395,0.9039622105855418,-0.38377548571655035,-0.9417824279857177,0.28491329175424573,0.9732271270498151,-0.17106684345077872,-0.9940766590333264,0.04285747872919846,0.999657726799591,0.09805152221776776,-0.985027376496916,-0.24868988716497914,
0.9452616647897091,0.4045472178879115,-0.8758624742544932,-0.5594135319425779,0.7732855634213638,0.7053456827732624,-0.6355765145327038,-0.8328192599541004,0.4630783014411666,0.9311267646590414,-0.2591453255417704,-0.9890740392187082,0.030766169093095375,0.9960041260451147,0.2110346319341552,-0.9431376225839149,
-0.4511699000511085,0.8251597619485228,0.670999860942617,-0.6419089236431357,-0.8495202811098108,0.39993625527105425,0.9653111125920658,-0.11362528897131971,-0.9992226935732867,-0.19449542546891307,0.9376240811868674,0.4946181638120598,-0.7758494632252803,-0.7519967101212217,0.521280465089589,0.9308801596315602,
-0.19533880186778324,-0.9998685450900215,-0.16640538080752737,0.9381355208580071,0.5167130042593379,-0.7415398935533003,-0.802139493349508,0.4272791970503417,0.9713317283040841,-0.03555422832648187,-0.9852594252640416,-0.3731444914245778,0.8276497743074627,0.7259343168357262,-0.5131854716652697,-0.9503709271486884,
0.09071413513929916,0.9905340690738222,0.3609182277571742,-0.8231770556884941,-0.7455646918621359,0.469598094501957,0.9700774057275657,0.001351222235442844,-0.9686747413782426,-0.48256080051416983,0.7253849404755924,0.8509751277300442,-0.28720854208608937,-0.9996447515291285,-0.2386825705196091,0.8719214500415734,
0.7070850658829174,-0.4870731199175568,-0.973886566865025,-0.05365461355310839,0.942953735405113,0.587636174758565,-0.6059191833873006,-0.9372391643801946,0.05837646291951751,0.9707742424068256,0.5193922790375888,-0.6577801294485379,-0.917888732123746,0.0951171842251602,0.9757758780563391,0.5136071276317543,
-0.6515122786401066,-0.9268998227344977,0.0568435329707618,0.9626986711387524,0.5711169734686521,-0.5859452362550388,-0.9593370929094306,-0.056720892737711526,0.9200201797783497,0.6827990092916144,-0.45045718935554424,-0.9936969735703642,-0.24315332620536376,0.8216046334379465,0.8251944560694946,-0.23116034784682868,
-0.9906684841625836,-0.48793114308331964,0.6327271278299522,0.9535305376404022,0.07590249324531644,-0.8956024966413276,-0.7506591446323682,0.32468723941967054,0.997991867054955,0.4443600886739411,-0.6520246743932532,-0.9531968580332627,-0.09878497455484683,0.8736900671497718,0.7957122431035348,-0.2333109866918325,
-0.9833638606885897,-0.5677847611442951,0.5165552417177618,0.9933197150904917,0.3093674522303538,-0.7332428174379773,-0.9260908906796308,-0.052305288699186166,0.880183576927755,0.8074255846108802,-0.18176747662315657,-0.9641796253014532,-0.6614270356027826,0.3809378743652582,0.9975882680365553,0.5079043511874277,
-0.5411057569891236,-0.9947568692207648,-0.3614909536531962,0.6635893314143555,0.9695833066135854,0.23193709834571716,-0.752846280056459,-0.9341186309057536,-0.12502855314728134,0.814611577151806,0.8979667705730853,0.043716541685519694,-0.8545359328173722,-0.8681975446019556,0.010809570652078056,0.8772813141294039,
0.8495202811096697,-0.038254831877669475,-0.8859758300466642,-0.8445253285208336,0.0386230747917501,0.8819266929427968,0.853865308257398,-0.01191504503112016,-0.8645167134414014,-0.8763066800439252,-0.041875653729171035,0.8312520164521842,0.9086343226759462,0.1224687749254994,-0.7779763094229916,-0.9454418975269331,
-0.2287096332866304,0.6993121972808145,0.9788945933977149,0.35770845281286356,-0.5894237869695266,-0.9986117983944375,-0.5037717663731474,0.443204251209147,0.991882081237177,0.6572711021616114,-0.2579587097435145,-0.9444773193549375,-0.8037137476363022,0.03555422832674925,0.8423475932975986,0.9234264326750142,
0.21517520593747957,-0.6744082097962316,-0.9923969604075246,-0.4762544056611531,0.43641960223758236,0.98486813025768,0.7194393454791972,-0.13556344345808757,-0.8781348357468007,-0.9072443241056106,-0.20526754444428627,0.6595362757447504,0.9973122276380169,0.5451282918804483,-0.33477644538895496,-0.9509425742390781,
-0.8268215661504691,-0.06450677023600318,0.7455237586507313,0.9850061919679485,0.477280202274066,-0.38876087467713627,-0.9616950233435587,-0.8178405810626352,-0.0697768969286048,0.7277060603809756,0.9920761651911643,0.5362934346887608,-0.3048082404095647,-0.9255569763537951,-0.8863173735938055,-0.22074985136408876,
0.5981215803145051,0.997626483190521,0.7046923159673673,-0.07265626914275577,-0.7982718948739636,-0.9796040563169521,-0.4993083629293127,0.3144443458494678,0.9166166325817039,0.9108780827064359,0.30673799752992364,-0.4958987477736227,-0.9749493844498841,-0.8251597619484309,-0.14833078149447007,0.6207626346405161,
0.9963474817979885,0.7471180684162626,0.034142444607836525,-0.6978619477542031,-0.9999866912863024,-0.6926084943183511,0.032423659700346656,0.7358683925902817,0.9988644148552395,0.6703164802777145,-0.050833189118322096,-0.7401785506422344,-0.9991176786215992,-0.6833373029149159,0.02112663674961348,0.7114579916888822,
0.9999304694126248,0.7298929372161397,0.05672089273789841,-0.6454811432944053,-0.9935376255187177,-0.8029090148808025,-0.18176747662362774,0.5342182281000675,0.9653912505854515,0.8886101900767628,0.3494354060781484,-0.36846716451062966,-0.8951101416022638,-0.9647799189938254,-0.5474432999270993,0.14249721801278203,
0.7593179370976132,0.999970055477208,0.7511458891695231,0.13909200518222956,-0.5376923700360762,-0.9556710295200649,-0.920140478427889,-0.45308730562146327,0.22308547290218372,0.7938858388287703,0.9993677485531182,0.7506591446324918,0.16513342248782012,-0.4918933579089748,-0.9288920324778026,-0.9568745665461746,
-0.568694473915292,0.06315830334384007,0.6656085971456042,0.9837741151906078,0.8875938723811243,0.4223306394684743,-0.21535514376757472,-0.7624663554937343,-0.9983970342055076,-0.8323770166568485,-0.33570228637772714,0.2913828346593136,0.8020294527387506,0.9999671357324733,0.8133628711426821,0.3182898011276006,
-0.29461263699280116,-0.7950049000991405,-0.9993936816673619,-0.8369436333696082,-0.37160543533355767,0.22524029545807567,0.7393520141142557,0.9906601112465891,0.8951101416023581,0.49060942465390367,-0.08000505513332462,-0.6209552261989727,-0.951113438890355,-0.9638039599022661,-0.6594439364759253,-0.14176767008864985,
0.4192104626939481,0.843833916364593,0.9999971311523869,0.8428768015140444,0.4257792915650769,-0.11966427385292795,-0.6262367667663898,-0.9426466165195914,-0.9779428121086001,-0.7261032626241473,-0.2647171523623591,0.27039842014603716,0.7260187952075616,0.9753304584204743,0.9523013511715133,0.6676230018007102,
0.2029226153782211,-0.3139195638370997,-0.7446225167480003,-0.9773617814374386,-0.9549083201156847,-0.687273428482953,-0.24654765490204353,0.25368368280895165,0.6882543272974337,0.9516808885117768,0.9830387597050245,0.778824563505633,0.39147540029074623,-0.08520783922224602,-0.5395036034244575,-0.8681060977762561,
-0.9991634991728605,-0.9070375492627036,-0.6160324660489052,-0.1929890389139486,0.2689198206150434,0.671136468750745,0.9306556045244146,0.996569527748079,0.8590961466716258,0.5497541260856779,0.13325069159264835,-0.30673799752972225,-0.68468141234178,-0.9296860181511639,-0.9982513437868271,-0.8811437714603633,
-0.6035222739865496,-0.2187725663864325,0.20238131206552637,0.5851984212256305,0.8641460441189653,0.9937313520640867,0.9552541427122613,0.7586380894609788,0.43940131858850034,0.05163059030603313,-0.3415968639976505,-0.678614680023552,-0.9086856122495266,-0.9992226935732899,-0.9397836161350681,-0.742486907165874,
-0.4390702548610516,-0.0752900586492556,0.2963142723637525,0.6241275672093204,0.8645167134410787,0.9873156684654814,0.9791199308720465,0.8441304078207613,0.6026404026684109,0.2875615115870699,-0.06039971911570213,-0.39819043769198026,-0.6857550264236422,-0.8906297874771946,-0.9913019737478629,-0.979044951334947,
-0.8581516320550341,-0.6446833125412893,-0.3640093246618578,-0.04752056609009044,0.27104880217977173,0.5592607933738403,0.7891941148339878,0.939951432649347,0.9992656645523431,0.9641307345666252,0.8404889618520441,0.6420972845792577,0.3887608746773312,0.10416195967636088,-0.1864762655696984,-0.458663198972474,
-0.6906566567090929,-0.8650718368290264,-0.9699878658803601,-0.999511371643157,-0.9538077137342182,-0.8386538419002695,-0.6645995709940413,-0.4458450789241147,-0.19895162854023468,0.058499091417478194,0.30919222855113876,0.5372262223597318,0.72905271060788,0.8741677155964148,0.9655352695373117,0.9997459657853027,
0.9769309469615577,0.9004657435602106,0.7765077985232477,0.6134164984892726,0.4211054495367702,0.21037418822073603,-0.007738743367515909,-0.22254659643730346,-0.42422259732337214,-0.6042076639800701,-0.7555081968643003,-0.8728821224020835,-0.9529179017251789,-0.9940164311586576,-0.9962895629968409,-0.9613913816528868,
-0.8922994824282162,-0.7930634806630179,-0.6685370293324389,-0.5241079628475387,-0.3654390341095832,-0.19822927778271263,-0.028003498983279817,0.1400650927990417,0.3012963886056101,0.45160834831227836,0.5875864778129374,0.7065202339836255,0.8064097983384665,0.8859473463574766,0.9444773193547266,0.9819403190726832,
0.9988051370273014,0.9959931481717528,0.9747988878636699,0.936810135545268,0.8838302863800558,0.8178052361511045,0.740756461745042,0.6547214702017018,0.5617023284573324,0.46362258320315747,0.36229254076522177,0.2593826018354532,0.15640413344736595,0.05469720669953626,-0.0445755723186253,-0.14042996583359413,
-0.2320565853100149,-0.3188137775677917,-0.40021770313477023,-0.4759303350785351,-0.5457460352564621,-0.6095772862509812,-0.6674400753625205,-0.7194393454790502,-0.7657548490340703,-0.8066276677020775,-0.8423475932974976,-0.8732415054398311,-0.8996628293427987,-0.9219821126250932,-0.9405787231433316,-0.9558336400523595,
-0.9681232870747527,-0.9778143396205302,-0.9852594252639776,-0.9907936294308151,-0.9947317142882849,-0.997365958116822,-0.9989645242676396,-0.9997702726522213,-0.9999999320982494,-0.9998435584446107,-0.9994642106138065,-0.9989977848253246,-0.9985529553977728,-0.9982111790780663,-0.9980267284283135,-0.9980267284283135);

end TestVectors;
